module johnson (input clk, output reg[3:0] = 4'b1000;
                always@(posedge clk)
                  begin
                    4'b0000:q=4'b1000;
                    4'b1000:q=4'b1100;
                    4'b1100:q=4'1110;
                    
