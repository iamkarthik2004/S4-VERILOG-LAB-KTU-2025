//Structureal flow
module possf(a,b,d,y)
  input a,b,d;
  output y;
  wire e,g,g;
  not (f,a,e);
  or (f,a,e);
  or(g,d,e);
endmodule
